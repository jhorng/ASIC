module Datapath_tb();

    reg Clock, Reset, IRload, JMPmux, PCload, Meminst, MemWr, Aload, Sub;
    reg [1:0]Asel;
    reg [7:0]Input;
    
    wire Aeq0, Apos;
    wire [7:5]IR;
    wire [7:0]Output, outputRam;
    wire [4:0]IR4_0, outputPC;
	
    integer i;

initial
begin
Clock=0;
Reset=1;
#2 Reset=0;
#2 start();
#2 fetch();
#2 decode();
#2 Input={$random}%256;
$display("value iDat!");
#2 load();
#2 inputState();
#2 writeMemory();
#2 add();
#10 sub();
#2 jz();
//#2 fetch();
//#2 decode();
#10 $finish;
end

initial
begin
$display("IRload | JMPmux | PCload | Meminst | MemWr | Aload | Sub |   Asel   |   Input  |  Output  |  outRam  |   IR   |  IR4_0  |  outputPC | time");
$monitor("	%b	%b	%b	%b	%b	%b	%b	%b	%b   %b   %b 	   %b 	   %b      %b %t", IRload, JMPmux, PCload, Meminst, MemWr, Aload, Sub, Asel, Input, Output, outputRam, IR, IR4_0, outputPC, $time);
end


task writeMemory;
begin
$display("Write data into memory!");
	for(i=0; i<3; i=i+1)
	begin
		#2 PCload=0;
		IRload=1;
		JMPmux=1;
		Meminst=0;
		MemWr=1;
		#2 Asel = 2'b01;
		Aload = 1;
		Input={$random}%256;
	end
	MemWr=0;
	Aload=0;
end
endtask

task oneTimeReset();
begin
$display("Clear register!");
  #2 Reset=1;
	IRload=0;
	JMPmux=0;
	PCload=0;
	Meminst=0;
	MemWr=0;
	Aload=0;
	Sub=0;
	Asel=0;
  #4 Reset=0;
end
endtask

task start;
begin
$display("Start!");
IRload=0;
JMPmux=0;
PCload=0;
Meminst=0;
MemWr=0;
Aload=0;
Sub=0;
Asel=0;
end
endtask

task fetch;
begin
$display("Fetch!");
IRload=1;
JMPmux=0;
PCload=1;
Meminst=0;
MemWr=0;
Aload=0;
Sub=0;
Asel=0;
end
endtask

task decode;
begin
$display("Decode!");
IRload=0;
JMPmux=0;
PCload=0;
Meminst=1;
MemWr=0;
Aload=0;
Sub=0;
Asel=0;
end
endtask

task load;
begin
$display("Load!");
IRload=0;
JMPmux=0;
PCload=0;
Meminst=0;
MemWr=0;
Aload=1;
Sub=0;
Asel=2'b10;
end
endtask

task store;
begin
$display("Store!");
IRload=0;
JMPmux=0;
PCload=0;
Meminst=1;
MemWr=1;
Aload=0;
Sub=0;
Asel=0;
end
endtask

task add;
begin
$display("Add!");
IRload=0;
JMPmux=0;
PCload=0;
Meminst=0;
MemWr=0;
Aload=1;
Sub=0;
Asel=0;
end
endtask

task sub;
begin
$display("Sub!");
IRload=0;
JMPmux=0;
PCload=0;
Meminst=0;
MemWr=0;
Aload=1;
Sub=1;
Asel=0;
end
endtask

task inputState;
begin
$display("Input!");
IRload=0;
JMPmux=0;
PCload=0;
Meminst=0;
MemWr=0;
Aload=1;
Sub=0;
Asel=2'b01;
Input={$random}%256;
end
endtask

task jz;
begin
$display("Jump if zero!");
IRload=0;
JMPmux=1;
PCload=Aeq0;
Meminst=0;
MemWr=0;
Aload=0;
Sub=0;
Asel=0;
end
endtask

task jpos;
begin
$display("Jump if positive!");
IRload=0;
JMPmux=1;
PCload=Apos;
Meminst=0;
MemWr=0;
Aload=0;
Sub=0;
Asel=0;
end
endtask

always #1 Clock=~Clock;

Datapath DP (Clock, Reset, IRload, JMPmux, PCload, Meminst, MemWr, Aload, Sub, Asel, Input, Aeq0, Apos, IR, Output, outputRam, IR4_0, outputPC);

endmodule 